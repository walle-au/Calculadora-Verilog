`timescale 1ns/1ps
// Sumador completo de 1 bit
module full_adder(
  input  wire a,
  input  wire b,
  input  wire cin,
  output wire sum,
  output wire cout
);
  assign {cout, sum} = a + b + cin;
endmodule
